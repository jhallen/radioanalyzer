module rom
  (
  clk,
  rd_addr,
  rd_data
  );

parameter ADDRWIDTH=8;
parameter WORDS = (1 << ADDRWIDTH);

input clk;

input [ADDRWIDTH-1:0] rd_addr;

output [31:0] rd_data;
reg [31:0] rd_data;

always @(posedge clk)
  case (rd_addr)
    16'h0000: rd_data <= 32'h00000093;
    16'h0001: rd_data <= 32'h00000193;
    16'h0002: rd_data <= 32'h00000213;
    16'h0003: rd_data <= 32'h00000293;
    16'h0004: rd_data <= 32'h00000313;
    16'h0005: rd_data <= 32'h00000393;
    16'h0006: rd_data <= 32'h00000413;
    16'h0007: rd_data <= 32'h00000493;
    16'h0008: rd_data <= 32'h00000513;
    16'h0009: rd_data <= 32'h00000593;
    16'h000a: rd_data <= 32'h00000613;
    16'h000b: rd_data <= 32'h00000693;
    16'h000c: rd_data <= 32'h00000713;
    16'h000d: rd_data <= 32'h00000793;
    16'h000e: rd_data <= 32'h00000813;
    16'h000f: rd_data <= 32'h00000893;
    16'h0010: rd_data <= 32'h00000913;
    16'h0011: rd_data <= 32'h00000993;
    16'h0012: rd_data <= 32'h00000a13;
    16'h0013: rd_data <= 32'h00000a93;
    16'h0014: rd_data <= 32'h00000b13;
    16'h0015: rd_data <= 32'h00000b93;
    16'h0016: rd_data <= 32'h00000c13;
    16'h0017: rd_data <= 32'h00000c93;
    16'h0018: rd_data <= 32'h00000d13;
    16'h0019: rd_data <= 32'h00000d93;
    16'h001a: rd_data <= 32'h00000e13;
    16'h001b: rd_data <= 32'h00000e93;
    16'h001c: rd_data <= 32'h00000f13;
    16'h001d: rd_data <= 32'h00000f93;
    16'h001e: rd_data <= 32'h03000537;
    16'h001f: rd_data <= 32'hc10c4585;
    16'h0020: rd_data <= 32'hc1084501;
    16'h0021: rd_data <= 32'h4ee30511;
    16'h0022: rd_data <= 32'h0537fe25;
    16'h0023: rd_data <= 32'h458d0300;
    16'h0024: rd_data <= 32'h2517c10c;
    16'h0025: rd_data <= 32'h05130000;
    16'h0026: rd_data <= 32'h0593a465;
    16'h0027: rd_data <= 32'h06130000;
    16'h0028: rd_data <= 32'hd8630000;
    16'h0029: rd_data <= 32'h411400c5;
    16'h002a: rd_data <= 32'h0511c194;
    16'h002b: rd_data <= 32'hcce30591;
    16'h002c: rd_data <= 32'h0537fec5;
    16'h002d: rd_data <= 32'h459d0300;
    16'h002e: rd_data <= 32'h0513c10c;
    16'h002f: rd_data <= 32'h05930000;
    16'h0030: rd_data <= 32'h57630000;
    16'h0031: rd_data <= 32'h202300b5;
    16'h0032: rd_data <= 32'h05110005;
    16'h0033: rd_data <= 32'hfeb54de3;
    16'h0034: rd_data <= 32'h03000537;
    16'h0035: rd_data <= 32'hc10c45bd;
    16'h0036: rd_data <= 32'h2a0010ef;
    16'h0037: rd_data <= 32'h0001a001;
    16'h0038: rd_data <= 32'h020002b7;
    16'h0039: rd_data <= 32'h12000313;
    16'h003a: rd_data <= 32'h00629023;
    16'h003b: rd_data <= 32'h000281a3;
    16'h003c: rd_data <= 32'h4f21c605;
    16'h003d: rd_data <= 32'h0ff67393;
    16'h003e: rd_data <= 32'h0073de93;
    16'h003f: rd_data <= 32'h01d28023;
    16'h0040: rd_data <= 32'h010eee93;
    16'h0041: rd_data <= 32'h01d28023;
    16'h0042: rd_data <= 32'hf3930386;
    16'h0043: rd_data <= 32'h1f7d0ff3;
    16'h0044: rd_data <= 32'hfe0f14e3;
    16'h0045: rd_data <= 32'h00628023;
    16'h0046: rd_data <= 32'h4f21cd9d;
    16'h0047: rd_data <= 32'h00054383;
    16'h0048: rd_data <= 32'h0073de93;
    16'h0049: rd_data <= 32'h01d28023;
    16'h004a: rd_data <= 32'h010eee93;
    16'h004b: rd_data <= 32'h01d28023;
    16'h004c: rd_data <= 32'h0002ce83;
    16'h004d: rd_data <= 32'h002efe93;
    16'h004e: rd_data <= 32'h001ede93;
    16'h004f: rd_data <= 32'he3b30386;
    16'h0050: rd_data <= 32'hf39301d3;
    16'h0051: rd_data <= 32'h1f7d0ff3;
    16'h0052: rd_data <= 32'hfc0f1ce3;
    16'h0053: rd_data <= 32'h00750023;
    16'h0054: rd_data <= 32'h15fd0505;
    16'h0055: rd_data <= 32'h0313b7d1;
    16'h0056: rd_data <= 32'h81a30800;
    16'h0057: rd_data <= 32'h80820062;
    16'h0058: rd_data <= 32'h71790000;
    16'h0059: rd_data <= 32'hd422d606;
    16'h005a: rd_data <= 32'h1800d226;
    16'h005b: rd_data <= 32'hfca42e23;
    16'h005c: rd_data <= 32'hfcb42c23;
    16'h005d: rd_data <= 32'hfcc40ba3;
    16'h005e: rd_data <= 32'h84b2860a;
    16'h005f: rd_data <= 32'h00010637;
    16'h0060: rd_data <= 32'h16060593;
    16'h0061: rd_data <= 32'h00010637;
    16'h0062: rd_data <= 32'h0e060613;
    16'h0063: rd_data <= 32'h40c58633;
    16'h0064: rd_data <= 32'h167d8609;
    16'h0065: rd_data <= 32'hfec42223;
    16'h0066: rd_data <= 32'h00010637;
    16'h0067: rd_data <= 32'h16060593;
    16'h0068: rd_data <= 32'h00010637;
    16'h0069: rd_data <= 32'h0e060613;
    16'h006a: rd_data <= 32'h40c58633;
    16'h006b: rd_data <= 32'h8e328609;
    16'h006c: rd_data <= 32'h56134e81;
    16'h006d: rd_data <= 32'h971301be;
    16'h006e: rd_data <= 32'h8f51005e;
    16'h006f: rd_data <= 32'h005e1693;
    16'h0070: rd_data <= 32'h00010737;
    16'h0071: rd_data <= 32'h16070693;
    16'h0072: rd_data <= 32'h00010737;
    16'h0073: rd_data <= 32'h0e070713;
    16'h0074: rd_data <= 32'h40e68733;
    16'h0075: rd_data <= 32'h833a8709;
    16'h0076: rd_data <= 32'h57134381;
    16'h0077: rd_data <= 32'h981301b3;
    16'h0078: rd_data <= 32'h68330053;
    16'h0079: rd_data <= 32'h17930107;
    16'h007a: rd_data <= 32'h07b70053;
    16'h007b: rd_data <= 32'h87130001;
    16'h007c: rd_data <= 32'h07b71607;
    16'h007d: rd_data <= 32'h87930001;
    16'h007e: rd_data <= 32'h07b30e07;
    16'h007f: rd_data <= 32'h078d40f7;
    16'h0080: rd_data <= 32'h07bd9bf1;
    16'h0081: rd_data <= 32'h07928391;
    16'h0082: rd_data <= 32'h40f10133;
    16'h0083: rd_data <= 32'h078d878a;
    16'h0084: rd_data <= 32'h078a8389;
    16'h0085: rd_data <= 32'hfef42023;
    16'h0086: rd_data <= 32'h000107b7;
    16'h0087: rd_data <= 32'h0e078793;
    16'h0088: rd_data <= 32'hfef42423;
    16'h0089: rd_data <= 32'hfe042783;
    16'h008a: rd_data <= 32'hfef42623;
    16'h008b: rd_data <= 32'h2703a839;
    16'h008c: rd_data <= 32'h0793fe84;
    16'h008d: rd_data <= 32'h24230047;
    16'h008e: rd_data <= 32'h2783fef4;
    16'h008f: rd_data <= 32'h8693fec4;
    16'h0090: rd_data <= 32'h26230047;
    16'h0091: rd_data <= 32'h4318fed4;
    16'h0092: rd_data <= 32'h2703c398;
    16'h0093: rd_data <= 32'h07b7fe84;
    16'h0094: rd_data <= 32'h87930001;
    16'h0095: rd_data <= 32'h1ce31607;
    16'h0096: rd_data <= 32'h2783fcf7;
    16'h0097: rd_data <= 32'h86befe04;
    16'h0098: rd_data <= 32'hfd842783;
    16'h0099: rd_data <= 32'hfd744703;
    16'h009a: rd_data <= 32'h85be863a;
    16'h009b: rd_data <= 32'hfdc42503;
    16'h009c: rd_data <= 32'h81269682;
    16'h009d: rd_data <= 32'h01130001;
    16'h009e: rd_data <= 32'h50b2fd04;
    16'h009f: rd_data <= 32'h54925422;
    16'h00a0: rd_data <= 32'h80826145;
    16'h00a1: rd_data <= 32'hce061101;
    16'h00a2: rd_data <= 32'h1000cc22;
    16'h00a3: rd_data <= 32'h008007b7;
    16'h00a4: rd_data <= 32'h26230789;
    16'h00a5: rd_data <= 32'h0793fef4;
    16'h00a6: rd_data <= 32'h00230650;
    16'h00a7: rd_data <= 32'h2783fef4;
    16'h00a8: rd_data <= 32'h83c1fec4;
    16'h00a9: rd_data <= 32'h0ff7f793;
    16'h00aa: rd_data <= 32'hfef400a3;
    16'h00ab: rd_data <= 32'hfec42783;
    16'h00ac: rd_data <= 32'hf79383a1;
    16'h00ad: rd_data <= 32'h01230ff7;
    16'h00ae: rd_data <= 32'h2783fef4;
    16'h00af: rd_data <= 32'hf793fec4;
    16'h00b0: rd_data <= 32'h01a30ff7;
    16'h00b1: rd_data <= 32'h0223fef4;
    16'h00b2: rd_data <= 32'h02a3fe04;
    16'h00b3: rd_data <= 32'h0793fe04;
    16'h00b4: rd_data <= 32'h4601fe04;
    16'h00b5: rd_data <= 32'h853e4599;
    16'h00b6: rd_data <= 32'h47833569;
    16'h00b7: rd_data <= 32'h05a3fe54;
    16'h00b8: rd_data <= 32'h0793fef4;
    16'h00b9: rd_data <= 32'h00230710;
    16'h00ba: rd_data <= 32'h2783fef4;
    16'h00bb: rd_data <= 32'h83c1fec4;
    16'h00bc: rd_data <= 32'h0ff7f793;
    16'h00bd: rd_data <= 32'hfef400a3;
    16'h00be: rd_data <= 32'hfec42783;
    16'h00bf: rd_data <= 32'hf79383a1;
    16'h00c0: rd_data <= 32'h01230ff7;
    16'h00c1: rd_data <= 32'h2783fef4;
    16'h00c2: rd_data <= 32'hf793fec4;
    16'h00c3: rd_data <= 32'h01a30ff7;
    16'h00c4: rd_data <= 32'h4783fef4;
    16'h00c5: rd_data <= 32'he793feb4;
    16'h00c6: rd_data <= 32'hf7930027;
    16'h00c7: rd_data <= 32'h02230ff7;
    16'h00c8: rd_data <= 32'h0793fef4;
    16'h00c9: rd_data <= 32'h4619fe04;
    16'h00ca: rd_data <= 32'h853e4595;
    16'h00cb: rd_data <= 32'h00013d1d;
    16'h00cc: rd_data <= 32'h446240f2;
    16'h00cd: rd_data <= 32'h80826105;
    16'h00ce: rd_data <= 32'hd6067179;
    16'h00cf: rd_data <= 32'h1800d422;
    16'h00d0: rd_data <= 32'h0fa387aa;
    16'h00d1: rd_data <= 32'h07b7fcf4;
    16'h00d2: rd_data <= 32'h43980200;
    16'h00d3: rd_data <= 32'hff8107b7;
    16'h00d4: rd_data <= 32'h76b317fd;
    16'h00d5: rd_data <= 32'h478300f7;
    16'h00d6: rd_data <= 32'h07c2fdf4;
    16'h00d7: rd_data <= 32'h07b7873e;
    16'h00d8: rd_data <= 32'h8f7d000f;
    16'h00d9: rd_data <= 32'h020007b7;
    16'h00da: rd_data <= 32'hc3988f55;
    16'h00db: rd_data <= 32'h008007b7;
    16'h00dc: rd_data <= 32'h26230791;
    16'h00dd: rd_data <= 32'h0793fef4;
    16'h00de: rd_data <= 32'h02230710;
    16'h00df: rd_data <= 32'h2783fef4;
    16'h00e0: rd_data <= 32'h83c1fec4;
    16'h00e1: rd_data <= 32'h0ff7f793;
    16'h00e2: rd_data <= 32'hfef402a3;
    16'h00e3: rd_data <= 32'hfec42783;
    16'h00e4: rd_data <= 32'hf79383a1;
    16'h00e5: rd_data <= 32'h03230ff7;
    16'h00e6: rd_data <= 32'h2783fef4;
    16'h00e7: rd_data <= 32'hf793fec4;
    16'h00e8: rd_data <= 32'h03a30ff7;
    16'h00e9: rd_data <= 32'h4783fef4;
    16'h00ea: rd_data <= 32'he793fdf4;
    16'h00eb: rd_data <= 32'hf7930707;
    16'h00ec: rd_data <= 32'h04230ff7;
    16'h00ed: rd_data <= 32'h0793fef4;
    16'h00ee: rd_data <= 32'h4619fe44;
    16'h00ef: rd_data <= 32'h853e4595;
    16'h00f0: rd_data <= 32'h0001334d;
    16'h00f1: rd_data <= 32'h542250b2;
    16'h00f2: rd_data <= 32'h80826145;
    16'h00f3: rd_data <= 32'hc6221141;
    16'h00f4: rd_data <= 32'h07b70800;
    16'h00f5: rd_data <= 32'h43940200;
    16'h00f6: rd_data <= 32'h020007b7;
    16'h00f7: rd_data <= 32'hff900737;
    16'h00f8: rd_data <= 32'h8f75177d;
    16'h00f9: rd_data <= 32'h0001c398;
    16'h00fa: rd_data <= 32'h01414432;
    16'h00fb: rd_data <= 32'h11418082;
    16'h00fc: rd_data <= 32'h0800c622;
    16'h00fd: rd_data <= 32'h020007b7;
    16'h00fe: rd_data <= 32'h07b74398;
    16'h00ff: rd_data <= 32'h17fdff90;
    16'h0100: rd_data <= 32'h00f776b3;
    16'h0101: rd_data <= 32'h020007b7;
    16'h0102: rd_data <= 32'h00400737;
    16'h0103: rd_data <= 32'hc3988f55;
    16'h0104: rd_data <= 32'h44320001;
    16'h0105: rd_data <= 32'h80820141;
    16'h0106: rd_data <= 32'hc6221141;
    16'h0107: rd_data <= 32'h07b70800;
    16'h0108: rd_data <= 32'h43980200;
    16'h0109: rd_data <= 32'hff9007b7;
    16'h010a: rd_data <= 32'h76b317fd;
    16'h010b: rd_data <= 32'h07b700f7;
    16'h010c: rd_data <= 32'h07370200;
    16'h010d: rd_data <= 32'h8f550020;
    16'h010e: rd_data <= 32'h0001c398;
    16'h010f: rd_data <= 32'h01414432;
    16'h0110: rd_data <= 32'h11418082;
    16'h0111: rd_data <= 32'h0800c622;
    16'h0112: rd_data <= 32'h020007b7;
    16'h0113: rd_data <= 32'h07b74398;
    16'h0114: rd_data <= 32'h17fdff90;
    16'h0115: rd_data <= 32'h00f776b3;
    16'h0116: rd_data <= 32'h020007b7;
    16'h0117: rd_data <= 32'h00600737;
    16'h0118: rd_data <= 32'hc3988f55;
    16'h0119: rd_data <= 32'h44320001;
    16'h011a: rd_data <= 32'h80820141;
    16'h011b: rd_data <= 32'hce061101;
    16'h011c: rd_data <= 32'h1000cc22;
    16'h011d: rd_data <= 32'h07a387aa;
    16'h011e: rd_data <= 32'h4703fef4;
    16'h011f: rd_data <= 32'h47a9fef4;
    16'h0120: rd_data <= 32'h00f71463;
    16'h0121: rd_data <= 32'h37dd4535;
    16'h0122: rd_data <= 32'h020007b7;
    16'h0123: rd_data <= 32'h470307a1;
    16'h0124: rd_data <= 32'hc398fef4;
    16'h0125: rd_data <= 32'h40f20001;
    16'h0126: rd_data <= 32'h61054462;
    16'h0127: rd_data <= 32'h11018082;
    16'h0128: rd_data <= 32'hcc22ce06;
    16'h0129: rd_data <= 32'h26231000;
    16'h012a: rd_data <= 32'ha819fea4;
    16'h012b: rd_data <= 32'hfec42783;
    16'h012c: rd_data <= 32'h00178713;
    16'h012d: rd_data <= 32'hfee42623;
    16'h012e: rd_data <= 32'h0007c783;
    16'h012f: rd_data <= 32'h377d853e;
    16'h0130: rd_data <= 32'hfec42783;
    16'h0131: rd_data <= 32'h0007c783;
    16'h0132: rd_data <= 32'h0001f3f5;
    16'h0133: rd_data <= 32'h446240f2;
    16'h0134: rd_data <= 32'h80826105;
    16'h0135: rd_data <= 32'hd6067179;
    16'h0136: rd_data <= 32'h1800d422;
    16'h0137: rd_data <= 32'hfca42e23;
    16'h0138: rd_data <= 32'hfcb42c23;
    16'h0139: rd_data <= 32'h2623479d;
    16'h013a: rd_data <= 32'ha8a9fef4;
    16'h013b: rd_data <= 32'hfec42783;
    16'h013c: rd_data <= 32'h2703078a;
    16'h013d: rd_data <= 32'h57b3fdc4;
    16'h013e: rd_data <= 32'hf71300f7;
    16'h013f: rd_data <= 32'h67c500f7;
    16'h0140: rd_data <= 32'h5c878793;
    16'h0141: rd_data <= 32'hc78397ba;
    16'h0142: rd_data <= 32'h05a30007;
    16'h0143: rd_data <= 32'h4703fef4;
    16'h0144: rd_data <= 32'h0793feb4;
    16'h0145: rd_data <= 32'h18630300;
    16'h0146: rd_data <= 32'h270300f7;
    16'h0147: rd_data <= 32'h2783fec4;
    16'h0148: rd_data <= 32'h5b63fd84;
    16'h0149: rd_data <= 32'h478300f7;
    16'h014a: rd_data <= 32'h853efeb4;
    16'h014b: rd_data <= 32'h27833781;
    16'h014c: rd_data <= 32'h2c23fec4;
    16'h014d: rd_data <= 32'ha011fcf4;
    16'h014e: rd_data <= 32'h27830001;
    16'h014f: rd_data <= 32'h17fdfec4;
    16'h0150: rd_data <= 32'hfef42623;
    16'h0151: rd_data <= 32'hfec42783;
    16'h0152: rd_data <= 32'hfa07d2e3;
    16'h0153: rd_data <= 32'h50b20001;
    16'h0154: rd_data <= 32'h61455422;
    16'h0155: rd_data <= 32'h11018082;
    16'h0156: rd_data <= 32'hcc22ce06;
    16'h0157: rd_data <= 32'h26231000;
    16'h0158: rd_data <= 32'h2703fea4;
    16'h0159: rd_data <= 32'h0793fec4;
    16'h015a: rd_data <= 32'hf7633e70;
    16'h015b: rd_data <= 32'h67c500e7;
    16'h015c: rd_data <= 32'h5dc78513;
    16'h015d: rd_data <= 32'hae05372d;
    16'h015e: rd_data <= 32'hfec42703;
    16'h015f: rd_data <= 32'h38300793;
    16'h0160: rd_data <= 32'h00e7fc63;
    16'h0161: rd_data <= 32'h03900513;
    16'h0162: rd_data <= 32'h278335d5;
    16'h0163: rd_data <= 32'h8793fec4;
    16'h0164: rd_data <= 32'h2623c7c7;
    16'h0165: rd_data <= 32'ha201fef4;
    16'h0166: rd_data <= 32'hfec42703;
    16'h0167: rd_data <= 32'h31f00793;
    16'h0168: rd_data <= 32'h00e7fc63;
    16'h0169: rd_data <= 32'h03800513;
    16'h016a: rd_data <= 32'h278335d1;
    16'h016b: rd_data <= 32'h8793fec4;
    16'h016c: rd_data <= 32'h2623ce07;
    16'h016d: rd_data <= 32'ha0c5fef4;
    16'h016e: rd_data <= 32'hfec42703;
    16'h016f: rd_data <= 32'h2bb00793;
    16'h0170: rd_data <= 32'h00e7fc63;
    16'h0171: rd_data <= 32'h03700513;
    16'h0172: rd_data <= 32'h27833555;
    16'h0173: rd_data <= 32'h8793fec4;
    16'h0174: rd_data <= 32'h2623d447;
    16'h0175: rd_data <= 32'ha0c1fef4;
    16'h0176: rd_data <= 32'hfec42703;
    16'h0177: rd_data <= 32'h25700793;
    16'h0178: rd_data <= 32'h00e7fc63;
    16'h0179: rd_data <= 32'h03600513;
    16'h017a: rd_data <= 32'h27833551;
    16'h017b: rd_data <= 32'h8793fec4;
    16'h017c: rd_data <= 32'h2623da87;
    16'h017d: rd_data <= 32'ha045fef4;
    16'h017e: rd_data <= 32'hfec42703;
    16'h017f: rd_data <= 32'h1f300793;
    16'h0180: rd_data <= 32'h00e7fc63;
    16'h0181: rd_data <= 32'h03500513;
    16'h0182: rd_data <= 32'h27833595;
    16'h0183: rd_data <= 32'h8793fec4;
    16'h0184: rd_data <= 32'h2623e0c7;
    16'h0185: rd_data <= 32'ha041fef4;
    16'h0186: rd_data <= 32'hfec42703;
    16'h0187: rd_data <= 32'h18f00793;
    16'h0188: rd_data <= 32'h00e7fc63;
    16'h0189: rd_data <= 32'h03400513;
    16'h018a: rd_data <= 32'h27833591;
    16'h018b: rd_data <= 32'h8793fec4;
    16'h018c: rd_data <= 32'h2623e707;
    16'h018d: rd_data <= 32'ha085fef4;
    16'h018e: rd_data <= 32'hfec42703;
    16'h018f: rd_data <= 32'h12b00793;
    16'h0190: rd_data <= 32'h00e7fc63;
    16'h0191: rd_data <= 32'h03300513;
    16'h0192: rd_data <= 32'h27833515;
    16'h0193: rd_data <= 32'h8793fec4;
    16'h0194: rd_data <= 32'h2623ed47;
    16'h0195: rd_data <= 32'ha081fef4;
    16'h0196: rd_data <= 32'hfec42703;
    16'h0197: rd_data <= 32'h0c700793;
    16'h0198: rd_data <= 32'h00e7fc63;
    16'h0199: rd_data <= 32'h03200513;
    16'h019a: rd_data <= 32'h27833511;
    16'h019b: rd_data <= 32'h8793fec4;
    16'h019c: rd_data <= 32'h2623f387;
    16'h019d: rd_data <= 32'ha005fef4;
    16'h019e: rd_data <= 32'hfec42703;
    16'h019f: rd_data <= 32'h06300793;
    16'h01a0: rd_data <= 32'h00e7fb63;
    16'h01a1: rd_data <= 32'h03100513;
    16'h01a2: rd_data <= 32'h278333d5;
    16'h01a3: rd_data <= 32'h8793fec4;
    16'h01a4: rd_data <= 32'h2623f9c7;
    16'h01a5: rd_data <= 32'h2703fef4;
    16'h01a6: rd_data <= 32'h0793fec4;
    16'h01a7: rd_data <= 32'hfc630590;
    16'h01a8: rd_data <= 32'h051300e7;
    16'h01a9: rd_data <= 32'h33d90390;
    16'h01aa: rd_data <= 32'hfec42783;
    16'h01ab: rd_data <= 32'hfa678793;
    16'h01ac: rd_data <= 32'hfef42623;
    16'h01ad: rd_data <= 32'h2703a8d5;
    16'h01ae: rd_data <= 32'h0793fec4;
    16'h01af: rd_data <= 32'hfc6304f0;
    16'h01b0: rd_data <= 32'h051300e7;
    16'h01b1: rd_data <= 32'h335d0380;
    16'h01b2: rd_data <= 32'hfec42783;
    16'h01b3: rd_data <= 32'hfb078793;
    16'h01b4: rd_data <= 32'hfef42623;
    16'h01b5: rd_data <= 32'h2703a8d1;
    16'h01b6: rd_data <= 32'h0793fec4;
    16'h01b7: rd_data <= 32'hfc630450;
    16'h01b8: rd_data <= 32'h051300e7;
    16'h01b9: rd_data <= 32'h33590370;
    16'h01ba: rd_data <= 32'hfec42783;
    16'h01bb: rd_data <= 32'hfba78793;
    16'h01bc: rd_data <= 32'hfef42623;
    16'h01bd: rd_data <= 32'h2703a855;
    16'h01be: rd_data <= 32'h0793fec4;
    16'h01bf: rd_data <= 32'hfc6303b0;
    16'h01c0: rd_data <= 32'h051300e7;
    16'h01c1: rd_data <= 32'h339d0360;
    16'h01c2: rd_data <= 32'hfec42783;
    16'h01c3: rd_data <= 32'hfc478793;
    16'h01c4: rd_data <= 32'hfef42623;
    16'h01c5: rd_data <= 32'h2703a851;
    16'h01c6: rd_data <= 32'h0793fec4;
    16'h01c7: rd_data <= 32'hfc630310;
    16'h01c8: rd_data <= 32'h051300e7;
    16'h01c9: rd_data <= 32'h33990350;
    16'h01ca: rd_data <= 32'hfec42783;
    16'h01cb: rd_data <= 32'hfce78793;
    16'h01cc: rd_data <= 32'hfef42623;
    16'h01cd: rd_data <= 32'h2703a895;
    16'h01ce: rd_data <= 32'h0793fec4;
    16'h01cf: rd_data <= 32'hfc630270;
    16'h01d0: rd_data <= 32'h051300e7;
    16'h01d1: rd_data <= 32'h331d0340;
    16'h01d2: rd_data <= 32'hfec42783;
    16'h01d3: rd_data <= 32'hfd878793;
    16'h01d4: rd_data <= 32'hfef42623;
    16'h01d5: rd_data <= 32'h2703a891;
    16'h01d6: rd_data <= 32'h47f5fec4;
    16'h01d7: rd_data <= 32'h00e7fb63;
    16'h01d8: rd_data <= 32'h03300513;
    16'h01d9: rd_data <= 32'h27833321;
    16'h01da: rd_data <= 32'h1789fec4;
    16'h01db: rd_data <= 32'hfef42623;
    16'h01dc: rd_data <= 32'h2703a825;
    16'h01dd: rd_data <= 32'h47cdfec4;
    16'h01de: rd_data <= 32'h00e7fb63;
    16'h01df: rd_data <= 32'h03200513;
    16'h01e0: rd_data <= 32'h278331f5;
    16'h01e1: rd_data <= 32'h17b1fec4;
    16'h01e2: rd_data <= 32'hfef42623;
    16'h01e3: rd_data <= 32'h2703a831;
    16'h01e4: rd_data <= 32'h47a5fec4;
    16'h01e5: rd_data <= 32'h00e7fa63;
    16'h01e6: rd_data <= 32'h03100513;
    16'h01e7: rd_data <= 32'h278339c1;
    16'h01e8: rd_data <= 32'h17d9fec4;
    16'h01e9: rd_data <= 32'hfef42623;
    16'h01ea: rd_data <= 32'hfec42703;
    16'h01eb: rd_data <= 32'hfb6347a1;
    16'h01ec: rd_data <= 32'h051300e7;
    16'h01ed: rd_data <= 32'h395d0390;
    16'h01ee: rd_data <= 32'hfec42783;
    16'h01ef: rd_data <= 32'h262317dd;
    16'h01f0: rd_data <= 32'ha0d5fef4;
    16'h01f1: rd_data <= 32'hfec42703;
    16'h01f2: rd_data <= 32'hfb63479d;
    16'h01f3: rd_data <= 32'h051300e7;
    16'h01f4: rd_data <= 32'h39690380;
    16'h01f5: rd_data <= 32'hfec42783;
    16'h01f6: rd_data <= 32'h262317e1;
    16'h01f7: rd_data <= 32'ha0e1fef4;
    16'h01f8: rd_data <= 32'hfec42703;
    16'h01f9: rd_data <= 32'hfb634799;
    16'h01fa: rd_data <= 32'h051300e7;
    16'h01fb: rd_data <= 32'h39bd0370;
    16'h01fc: rd_data <= 32'hfec42783;
    16'h01fd: rd_data <= 32'h262317e5;
    16'h01fe: rd_data <= 32'ha075fef4;
    16'h01ff: rd_data <= 32'hfec42703;
    16'h0200: rd_data <= 32'hfb634795;
    16'h0201: rd_data <= 32'h051300e7;
    16'h0202: rd_data <= 32'h318d0360;
    16'h0203: rd_data <= 32'hfec42783;
    16'h0204: rd_data <= 32'h262317e9;
    16'h0205: rd_data <= 32'ha841fef4;
    16'h0206: rd_data <= 32'hfec42703;
    16'h0207: rd_data <= 32'hfb634791;
    16'h0208: rd_data <= 32'h051300e7;
    16'h0209: rd_data <= 32'h31990350;
    16'h020a: rd_data <= 32'hfec42783;
    16'h020b: rd_data <= 32'h262317ed;
    16'h020c: rd_data <= 32'ha895fef4;
    16'h020d: rd_data <= 32'hfec42703;
    16'h020e: rd_data <= 32'hfb63478d;
    16'h020f: rd_data <= 32'h051300e7;
    16'h0210: rd_data <= 32'h312d0340;
    16'h0211: rd_data <= 32'hfec42783;
    16'h0212: rd_data <= 32'h262317f1;
    16'h0213: rd_data <= 32'ha8a1fef4;
    16'h0214: rd_data <= 32'hfec42703;
    16'h0215: rd_data <= 32'hfb634789;
    16'h0216: rd_data <= 32'h051300e7;
    16'h0217: rd_data <= 32'h31390330;
    16'h0218: rd_data <= 32'hfec42783;
    16'h0219: rd_data <= 32'h262317f5;
    16'h021a: rd_data <= 32'ha835fef4;
    16'h021b: rd_data <= 32'hfec42703;
    16'h021c: rd_data <= 32'hfb634785;
    16'h021d: rd_data <= 32'h051300e7;
    16'h021e: rd_data <= 32'h3ecd0320;
    16'h021f: rd_data <= 32'hfec42783;
    16'h0220: rd_data <= 32'h262317f9;
    16'h0221: rd_data <= 32'ha005fef4;
    16'h0222: rd_data <= 32'hfec42783;
    16'h0223: rd_data <= 32'h0513cb91;
    16'h0224: rd_data <= 32'h3ee90310;
    16'h0225: rd_data <= 32'hfec42783;
    16'h0226: rd_data <= 32'h262317fd;
    16'h0227: rd_data <= 32'ha021fef4;
    16'h0228: rd_data <= 32'h03000513;
    16'h0229: rd_data <= 32'h40f236e1;
    16'h022a: rd_data <= 32'h61054462;
    16'h022b: rd_data <= 32'h71798082;
    16'h022c: rd_data <= 32'hd422d606;
    16'h022d: rd_data <= 32'h2e231800;
    16'h022e: rd_data <= 32'h57fdfca4;
    16'h022f: rd_data <= 32'hfef42623;
    16'h0230: rd_data <= 32'hc00027f3;
    16'h0231: rd_data <= 32'hfef42423;
    16'h0232: rd_data <= 32'h030007b7;
    16'h0233: rd_data <= 32'hc398577d;
    16'h0234: rd_data <= 32'hfdc42783;
    16'h0235: rd_data <= 32'h2503c3ad;
    16'h0236: rd_data <= 32'h36d1fdc4;
    16'h0237: rd_data <= 32'h27f3a8a9;
    16'h0238: rd_data <= 32'h2223c000;
    16'h0239: rd_data <= 32'h2703fef4;
    16'h023a: rd_data <= 32'h2783fe44;
    16'h023b: rd_data <= 32'h07b3fe84;
    16'h023c: rd_data <= 32'h202340f7;
    16'h023d: rd_data <= 32'h2703fef4;
    16'h023e: rd_data <= 32'h27b7fe04;
    16'h023f: rd_data <= 32'h879300b7;
    16'h0240: rd_data <= 32'hf463b007;
    16'h0241: rd_data <= 32'h278302e7;
    16'h0242: rd_data <= 32'hc781fdc4;
    16'h0243: rd_data <= 32'hfdc42503;
    16'h0244: rd_data <= 32'h27833679;
    16'h0245: rd_data <= 32'h2423fe44;
    16'h0246: rd_data <= 32'h07b7fef4;
    16'h0247: rd_data <= 32'h43980300;
    16'h0248: rd_data <= 32'h030007b7;
    16'h0249: rd_data <= 32'hfff74713;
    16'h024a: rd_data <= 32'h07b7c398;
    16'h024b: rd_data <= 32'h07a10200;
    16'h024c: rd_data <= 32'h2623439c;
    16'h024d: rd_data <= 32'h2703fef4;
    16'h024e: rd_data <= 32'h57fdfec4;
    16'h024f: rd_data <= 32'hfaf701e3;
    16'h0250: rd_data <= 32'h030007b7;
    16'h0251: rd_data <= 32'h0007a023;
    16'h0252: rd_data <= 32'hfec42783;
    16'h0253: rd_data <= 32'h0ff7f793;
    16'h0254: rd_data <= 32'h50b2853e;
    16'h0255: rd_data <= 32'h61455422;
    16'h0256: rd_data <= 32'h11418082;
    16'h0257: rd_data <= 32'hc422c606;
    16'h0258: rd_data <= 32'h45010800;
    16'h0259: rd_data <= 32'h87aa37a9;
    16'h025a: rd_data <= 32'h40b2853e;
    16'h025b: rd_data <= 32'h01414422;
    16'h025c: rd_data <= 32'h11418082;
    16'h025d: rd_data <= 32'hc422c606;
    16'h025e: rd_data <= 32'h67c50800;
    16'h025f: rd_data <= 32'h5e478513;
    16'h0260: rd_data <= 32'h67c53e39;
    16'h0261: rd_data <= 32'h5f078513;
    16'h0262: rd_data <= 32'h07b73e19;
    16'h0263: rd_data <= 32'h439c0200;
    16'h0264: rd_data <= 32'h8bbd83c1;
    16'h0265: rd_data <= 32'h36c1853e;
    16'h0266: rd_data <= 32'h851367c5;
    16'h0267: rd_data <= 32'h36015fc7;
    16'h0268: rd_data <= 32'h851367c5;
    16'h0269: rd_data <= 32'h3ce56007;
    16'h026a: rd_data <= 32'h020007b7;
    16'h026b: rd_data <= 32'h07b74398;
    16'h026c: rd_data <= 32'h8ff90040;
    16'h026d: rd_data <= 32'h67c5c791;
    16'h026e: rd_data <= 32'h60878513;
    16'h026f: rd_data <= 32'ha02934cd;
    16'h0270: rd_data <= 32'h851367c5;
    16'h0271: rd_data <= 32'h3ce160c7;
    16'h0272: rd_data <= 32'h851367c5;
    16'h0273: rd_data <= 32'h3cc16147;
    16'h0274: rd_data <= 32'h020007b7;
    16'h0275: rd_data <= 32'h07b74398;
    16'h0276: rd_data <= 32'h8ff90020;
    16'h0277: rd_data <= 32'h67c5c791;
    16'h0278: rd_data <= 32'h60878513;
    16'h0279: rd_data <= 32'ha0293c6d;
    16'h027a: rd_data <= 32'h851367c5;
    16'h027b: rd_data <= 32'h3c4560c7;
    16'h027c: rd_data <= 32'h851367c5;
    16'h027d: rd_data <= 32'h346561c7;
    16'h027e: rd_data <= 32'h020007b7;
    16'h027f: rd_data <= 32'h07b74398;
    16'h0280: rd_data <= 32'h8ff90010;
    16'h0281: rd_data <= 32'h67c5c791;
    16'h0282: rd_data <= 32'h60878513;
    16'h0283: rd_data <= 32'ha0293c49;
    16'h0284: rd_data <= 32'h851367c5;
    16'h0285: rd_data <= 32'h346160c7;
    16'h0286: rd_data <= 32'h40b20001;
    16'h0287: rd_data <= 32'h01414422;
    16'h0288: rd_data <= 32'h71798082;
    16'h0289: rd_data <= 32'h1800d622;
    16'h028a: rd_data <= 32'hfca42e23;
    16'h028b: rd_data <= 32'hfdc42783;
    16'h028c: rd_data <= 32'h2623439c;
    16'h028d: rd_data <= 32'h2783fef4;
    16'h028e: rd_data <= 32'h07b6fec4;
    16'h028f: rd_data <= 32'hfec42703;
    16'h0290: rd_data <= 32'h26238fb9;
    16'h0291: rd_data <= 32'h2783fef4;
    16'h0292: rd_data <= 32'h83c5fec4;
    16'h0293: rd_data <= 32'hfec42703;
    16'h0294: rd_data <= 32'h26238fb9;
    16'h0295: rd_data <= 32'h2783fef4;
    16'h0296: rd_data <= 32'h0796fec4;
    16'h0297: rd_data <= 32'hfec42703;
    16'h0298: rd_data <= 32'h26238fb9;
    16'h0299: rd_data <= 32'h2783fef4;
    16'h029a: rd_data <= 32'h2703fdc4;
    16'h029b: rd_data <= 32'hc398fec4;
    16'h029c: rd_data <= 32'hfec42783;
    16'h029d: rd_data <= 32'h5432853e;
    16'h029e: rd_data <= 32'h80826145;
    16'h029f: rd_data <= 32'hde067139;
    16'h02a0: rd_data <= 32'hda26dc22;
    16'h02a1: rd_data <= 32'h47950080;
    16'h02a2: rd_data <= 32'hfcf42c23;
    16'h02a3: rd_data <= 32'h10000793;
    16'h02a4: rd_data <= 32'hfcf42a23;
    16'h02a5: rd_data <= 32'hfc042823;
    16'h02a6: rd_data <= 32'hfc042623;
    16'h02a7: rd_data <= 32'h851367c5;
    16'h02a8: rd_data <= 32'h3af56247;
    16'h02a9: rd_data <= 32'h26234785;
    16'h02aa: rd_data <= 32'ha855fef4;
    16'h02ab: rd_data <= 32'hfec42783;
    16'h02ac: rd_data <= 32'hfcf42423;
    16'h02ad: rd_data <= 32'hfe042423;
    16'h02ae: rd_data <= 32'h2783a02d;
    16'h02af: rd_data <= 32'h078afe84;
    16'h02b0: rd_data <= 32'hfd042703;
    16'h02b1: rd_data <= 32'h00f704b3;
    16'h02b2: rd_data <= 32'hfc840793;
    16'h02b3: rd_data <= 32'h3f91853e;
    16'h02b4: rd_data <= 32'hc09c87aa;
    16'h02b5: rd_data <= 32'hfe842703;
    16'h02b6: rd_data <= 32'hfd442783;
    16'h02b7: rd_data <= 32'h242397ba;
    16'h02b8: rd_data <= 32'h2703fef4;
    16'h02b9: rd_data <= 32'h67a1fe84;
    16'h02ba: rd_data <= 32'hfcf769e3;
    16'h02bb: rd_data <= 32'hfec42783;
    16'h02bc: rd_data <= 32'hfcf42423;
    16'h02bd: rd_data <= 32'hfe042223;
    16'h02be: rd_data <= 32'h2783a0a9;
    16'h02bf: rd_data <= 32'h078afe44;
    16'h02c0: rd_data <= 32'hfd042703;
    16'h02c1: rd_data <= 32'h438497ba;
    16'h02c2: rd_data <= 32'hfc840793;
    16'h02c3: rd_data <= 32'h3f11853e;
    16'h02c4: rd_data <= 32'h816387aa;
    16'h02c5: rd_data <= 32'h67c502f4;
    16'h02c6: rd_data <= 32'h63878513;
    16'h02c7: rd_data <= 32'h27833249;
    16'h02c8: rd_data <= 32'h078afe44;
    16'h02c9: rd_data <= 32'h853e4591;
    16'h02ca: rd_data <= 32'h67c53275;
    16'h02cb: rd_data <= 32'h5fc78513;
    16'h02cc: rd_data <= 32'ha0e132bd;
    16'h02cd: rd_data <= 32'hfe442703;
    16'h02ce: rd_data <= 32'hfd442783;
    16'h02cf: rd_data <= 32'h222397ba;
    16'h02d0: rd_data <= 32'h2703fef4;
    16'h02d1: rd_data <= 32'h67a1fe44;
    16'h02d2: rd_data <= 32'hfaf769e3;
    16'h02d3: rd_data <= 32'h851367c5;
    16'h02d4: rd_data <= 32'h32b16507;
    16'h02d5: rd_data <= 32'hfec42783;
    16'h02d6: rd_data <= 32'h26230785;
    16'h02d7: rd_data <= 32'h2703fef4;
    16'h02d8: rd_data <= 32'h2783fec4;
    16'h02d9: rd_data <= 32'hd3e3fd84;
    16'h02da: rd_data <= 32'h2023f4e7;
    16'h02db: rd_data <= 32'ha00dfe04;
    16'h02dc: rd_data <= 32'hfe042783;
    16'h02dd: rd_data <= 32'hfcc42703;
    16'h02de: rd_data <= 32'h270397ba;
    16'h02df: rd_data <= 32'h7713fe04;
    16'h02e0: rd_data <= 32'h80230ff7;
    16'h02e1: rd_data <= 32'h278300e7;
    16'h02e2: rd_data <= 32'h0785fe04;
    16'h02e3: rd_data <= 32'hfef42023;
    16'h02e4: rd_data <= 32'hfe042703;
    16'h02e5: rd_data <= 32'h07f00793;
    16'h02e6: rd_data <= 32'hfce7dce3;
    16'h02e7: rd_data <= 32'hfc042e23;
    16'h02e8: rd_data <= 32'h2783a099;
    16'h02e9: rd_data <= 32'h2703fdc4;
    16'h02ea: rd_data <= 32'h97bafcc4;
    16'h02eb: rd_data <= 32'h0007c783;
    16'h02ec: rd_data <= 32'h0ff7f713;
    16'h02ed: rd_data <= 32'hfdc42783;
    16'h02ee: rd_data <= 32'h0ff7f793;
    16'h02ef: rd_data <= 32'h02f70063;
    16'h02f0: rd_data <= 32'h851367c5;
    16'h02f1: rd_data <= 32'h38e16547;
    16'h02f2: rd_data <= 32'hfdc42783;
    16'h02f3: rd_data <= 32'h853e4591;
    16'h02f4: rd_data <= 32'h67c53211;
    16'h02f5: rd_data <= 32'h5fc78513;
    16'h02f6: rd_data <= 32'ha00530d9;
    16'h02f7: rd_data <= 32'hfdc42783;
    16'h02f8: rd_data <= 32'h2e230785;
    16'h02f9: rd_data <= 32'h2703fcf4;
    16'h02fa: rd_data <= 32'h0793fdc4;
    16'h02fb: rd_data <= 32'hdae307f0;
    16'h02fc: rd_data <= 32'h67c5fae7;
    16'h02fd: rd_data <= 32'h66c78513;
    16'h02fe: rd_data <= 32'h50f2305d;
    16'h02ff: rd_data <= 32'h54d25462;
    16'h0300: rd_data <= 32'h80826121;
    16'h0301: rd_data <= 32'hd6067179;
    16'h0302: rd_data <= 32'h1800d422;
    16'h0303: rd_data <= 32'hfc042c23;
    16'h0304: rd_data <= 32'hfc042e23;
    16'h0305: rd_data <= 32'hfe042023;
    16'h0306: rd_data <= 32'hfe042223;
    16'h0307: rd_data <= 32'hfe040423;
    16'h0308: rd_data <= 32'hf9f00793;
    16'h0309: rd_data <= 32'hfcf40c23;
    16'h030a: rd_data <= 32'hfd840793;
    16'h030b: rd_data <= 32'h45c54601;
    16'h030c: rd_data <= 32'hf0ef853e;
    16'h030d: rd_data <= 32'h4785d30f;
    16'h030e: rd_data <= 32'hfef42623;
    16'h030f: rd_data <= 32'h0513a01d;
    16'h0310: rd_data <= 32'h302d0200;
    16'h0311: rd_data <= 32'hfec42783;
    16'h0312: rd_data <= 32'hff040713;
    16'h0313: rd_data <= 32'hc78397ba;
    16'h0314: rd_data <= 32'h4589fe87;
    16'h0315: rd_data <= 32'h38bd853e;
    16'h0316: rd_data <= 32'hfec42783;
    16'h0317: rd_data <= 32'h26230785;
    16'h0318: rd_data <= 32'h2703fef4;
    16'h0319: rd_data <= 32'h47c1fec4;
    16'h031a: rd_data <= 32'hfce7dbe3;
    16'h031b: rd_data <= 32'hf0ef4529;
    16'h031c: rd_data <= 32'h0001ffef;
    16'h031d: rd_data <= 32'h542250b2;
    16'h031e: rd_data <= 32'h80826145;
    16'h031f: rd_data <= 32'hd6067179;
    16'h0320: rd_data <= 32'h1800d422;
    16'h0321: rd_data <= 32'hfca42e23;
    16'h0322: rd_data <= 32'hfcb42c23;
    16'h0323: rd_data <= 32'hf0ef4521;
    16'h0324: rd_data <= 32'h0793eaaf;
    16'h0325: rd_data <= 32'h04230650;
    16'h0326: rd_data <= 32'h2783fef4;
    16'h0327: rd_data <= 32'h83c1fdc4;
    16'h0328: rd_data <= 32'h0ff7f793;
    16'h0329: rd_data <= 32'hfef404a3;
    16'h032a: rd_data <= 32'hfdc42783;
    16'h032b: rd_data <= 32'hf79383a1;
    16'h032c: rd_data <= 32'h05230ff7;
    16'h032d: rd_data <= 32'h2783fef4;
    16'h032e: rd_data <= 32'hf793fdc4;
    16'h032f: rd_data <= 32'h05a30ff7;
    16'h0330: rd_data <= 32'h0623fef4;
    16'h0331: rd_data <= 32'h06a3fe04;
    16'h0332: rd_data <= 32'h0793fe04;
    16'h0333: rd_data <= 32'h4601fe84;
    16'h0334: rd_data <= 32'h853e4599;
    16'h0335: rd_data <= 32'hc8eff0ef;
    16'h0336: rd_data <= 32'h851367c5;
    16'h0337: rd_data <= 32'hf0ef6787;
    16'h0338: rd_data <= 32'h4599fc0f;
    16'h0339: rd_data <= 32'hfdc42503;
    16'h033a: rd_data <= 32'hfecff0ef;
    16'h033b: rd_data <= 32'h851367c5;
    16'h033c: rd_data <= 32'hf0ef67c7;
    16'h033d: rd_data <= 32'h2503facf;
    16'h033e: rd_data <= 32'hf0effd84;
    16'h033f: rd_data <= 32'h67c5fa4f;
    16'h0340: rd_data <= 32'h68078513;
    16'h0341: rd_data <= 32'hf9aff0ef;
    16'h0342: rd_data <= 32'hfed44783;
    16'h0343: rd_data <= 32'h853e4589;
    16'h0344: rd_data <= 32'hfc4ff0ef;
    16'h0345: rd_data <= 32'h851367c5;
    16'h0346: rd_data <= 32'hf0ef5fc7;
    16'h0347: rd_data <= 32'h4783f84f;
    16'h0348: rd_data <= 32'h853efed4;
    16'h0349: rd_data <= 32'h542250b2;
    16'h034a: rd_data <= 32'h80826145;
    16'h034b: rd_data <= 32'hce061101;
    16'h034c: rd_data <= 32'h1000cc22;
    16'h034d: rd_data <= 32'h851367c5;
    16'h034e: rd_data <= 32'hf0ef5fc7;
    16'h034f: rd_data <= 32'h67c5f64f;
    16'h0350: rd_data <= 32'h68478593;
    16'h0351: rd_data <= 32'h00800537;
    16'h0352: rd_data <= 32'h87aa3f15;
    16'h0353: rd_data <= 32'hfef407a3;
    16'h0354: rd_data <= 32'h859367c5;
    16'h0355: rd_data <= 32'h07b768c7;
    16'h0356: rd_data <= 32'h85130080;
    16'h0357: rd_data <= 32'h3f390017;
    16'h0358: rd_data <= 32'h072387aa;
    16'h0359: rd_data <= 32'h67c5fef4;
    16'h035a: rd_data <= 32'h69478593;
    16'h035b: rd_data <= 32'h008007b7;
    16'h035c: rd_data <= 32'h00278513;
    16'h035d: rd_data <= 32'h87aa3721;
    16'h035e: rd_data <= 32'hfef406a3;
    16'h035f: rd_data <= 32'h859367c5;
    16'h0360: rd_data <= 32'h07b769c7;
    16'h0361: rd_data <= 32'h85130080;
    16'h0362: rd_data <= 32'h3dcd0037;
    16'h0363: rd_data <= 32'h062387aa;
    16'h0364: rd_data <= 32'h67c5fef4;
    16'h0365: rd_data <= 32'h6a478593;
    16'h0366: rd_data <= 32'h008007b7;
    16'h0367: rd_data <= 32'h00478513;
    16'h0368: rd_data <= 32'h87aa3df1;
    16'h0369: rd_data <= 32'hfef405a3;
    16'h036a: rd_data <= 32'h859367c5;
    16'h036b: rd_data <= 32'h07b76ac7;
    16'h036c: rd_data <= 32'h85130080;
    16'h036d: rd_data <= 32'h35d90057;
    16'h036e: rd_data <= 32'h052387aa;
    16'h036f: rd_data <= 32'h0001fef4;
    16'h0370: rd_data <= 32'h446240f2;
    16'h0371: rd_data <= 32'h80826105;
    16'h0372: rd_data <= 32'h2623714d;
    16'h0373: rd_data <= 32'h24231411;
    16'h0374: rd_data <= 32'h0a801481;
    16'h0375: rd_data <= 32'h2c2387aa;
    16'h0376: rd_data <= 32'h0fa3eab4;
    16'h0377: rd_data <= 32'h0793eaf4;
    16'h0378: rd_data <= 32'h2a23ec04;
    16'h0379: rd_data <= 32'hb7b7fcf4;
    16'h037a: rd_data <= 32'h879312b9;
    16'h037b: rd_data <= 32'h26230a17;
    16'h037c: rd_data <= 32'h27f3fef4;
    16'h037d: rd_data <= 32'h2823c000;
    16'h037e: rd_data <= 32'h27f3fcf4;
    16'h037f: rd_data <= 32'h2623c020;
    16'h0380: rd_data <= 32'h2423fcf4;
    16'h0381: rd_data <= 32'ha8d5fe04;
    16'h0382: rd_data <= 32'hfe042223;
    16'h0383: rd_data <= 32'h2783a889;
    16'h0384: rd_data <= 32'h07b6fec4;
    16'h0385: rd_data <= 32'hfec42703;
    16'h0386: rd_data <= 32'h26238fb9;
    16'h0387: rd_data <= 32'h2783fef4;
    16'h0388: rd_data <= 32'h83c5fec4;
    16'h0389: rd_data <= 32'hfec42703;
    16'h038a: rd_data <= 32'h26238fb9;
    16'h038b: rd_data <= 32'h2783fef4;
    16'h038c: rd_data <= 32'h0796fec4;
    16'h038d: rd_data <= 32'hfec42703;
    16'h038e: rd_data <= 32'h26238fb9;
    16'h038f: rd_data <= 32'h2783fef4;
    16'h0390: rd_data <= 32'hf713fec4;
    16'h0391: rd_data <= 32'h27830ff7;
    16'h0392: rd_data <= 32'h0693fe44;
    16'h0393: rd_data <= 32'h97b6ff04;
    16'h0394: rd_data <= 32'hece78823;
    16'h0395: rd_data <= 32'hfe442783;
    16'h0396: rd_data <= 32'h22230785;
    16'h0397: rd_data <= 32'h2703fef4;
    16'h0398: rd_data <= 32'h0793fe44;
    16'h0399: rd_data <= 32'hd4e30ff0;
    16'h039a: rd_data <= 32'h2023fae7;
    16'h039b: rd_data <= 32'h2e23fe04;
    16'h039c: rd_data <= 32'ha82dfc04;
    16'h039d: rd_data <= 32'hfe042783;
    16'h039e: rd_data <= 32'hff040713;
    16'h039f: rd_data <= 32'hc78397ba;
    16'h03a0: rd_data <= 32'hc385ed07;
    16'h03a1: rd_data <= 32'hfdc42783;
    16'h03a2: rd_data <= 32'h00178713;
    16'h03a3: rd_data <= 32'hfce42e23;
    16'h03a4: rd_data <= 32'hfe042703;
    16'h03a5: rd_data <= 32'h0ff77713;
    16'h03a6: rd_data <= 32'hff040693;
    16'h03a7: rd_data <= 32'h882397b6;
    16'h03a8: rd_data <= 32'h2783ece7;
    16'h03a9: rd_data <= 32'h0785fe04;
    16'h03aa: rd_data <= 32'hfef42023;
    16'h03ab: rd_data <= 32'hfe042703;
    16'h03ac: rd_data <= 32'h0ff00793;
    16'h03ad: rd_data <= 32'hfce7d0e3;
    16'h03ae: rd_data <= 32'hfc042c23;
    16'h03af: rd_data <= 32'hfc042423;
    16'h03b0: rd_data <= 32'h2783a015;
    16'h03b1: rd_data <= 32'h078afd84;
    16'h03b2: rd_data <= 32'hfd442703;
    16'h03b3: rd_data <= 32'h439c97ba;
    16'h03b4: rd_data <= 32'hfec42703;
    16'h03b5: rd_data <= 32'h26238fb9;
    16'h03b6: rd_data <= 32'h2783fef4;
    16'h03b7: rd_data <= 32'h0785fd84;
    16'h03b8: rd_data <= 32'hfcf42c23;
    16'h03b9: rd_data <= 32'hfd842703;
    16'h03ba: rd_data <= 32'h03f00793;
    16'h03bb: rd_data <= 32'hfce7dbe3;
    16'h03bc: rd_data <= 32'hfe842783;
    16'h03bd: rd_data <= 32'h24230785;
    16'h03be: rd_data <= 32'h2703fef4;
    16'h03bf: rd_data <= 32'h47cdfe84;
    16'h03c0: rd_data <= 32'hf0e7d4e3;
    16'h03c1: rd_data <= 32'hc00027f3;
    16'h03c2: rd_data <= 32'hfcf42223;
    16'h03c3: rd_data <= 32'hc02027f3;
    16'h03c4: rd_data <= 32'hfcf42023;
    16'h03c5: rd_data <= 32'hebf44783;
    16'h03c6: rd_data <= 32'h67c5c3b5;
    16'h03c7: rd_data <= 32'h6b478513;
    16'h03c8: rd_data <= 32'hd7eff0ef;
    16'h03c9: rd_data <= 32'hfc442703;
    16'h03ca: rd_data <= 32'hfd042783;
    16'h03cb: rd_data <= 32'h40f707b3;
    16'h03cc: rd_data <= 32'h853e45a1;
    16'h03cd: rd_data <= 32'hda0ff0ef;
    16'h03ce: rd_data <= 32'hf0ef4529;
    16'h03cf: rd_data <= 32'h67c5d32f;
    16'h03d0: rd_data <= 32'h6c078513;
    16'h03d1: rd_data <= 32'hd5aff0ef;
    16'h03d2: rd_data <= 32'hfc042703;
    16'h03d3: rd_data <= 32'hfcc42783;
    16'h03d4: rd_data <= 32'h40f707b3;
    16'h03d5: rd_data <= 32'h853e45a1;
    16'h03d6: rd_data <= 32'hd7cff0ef;
    16'h03d7: rd_data <= 32'hf0ef4529;
    16'h03d8: rd_data <= 32'h67c5d0ef;
    16'h03d9: rd_data <= 32'h6cc78513;
    16'h03da: rd_data <= 32'hd36ff0ef;
    16'h03db: rd_data <= 32'h250345a1;
    16'h03dc: rd_data <= 32'hf0effec4;
    16'h03dd: rd_data <= 32'h4529d62f;
    16'h03de: rd_data <= 32'hcf4ff0ef;
    16'h03df: rd_data <= 32'heb842783;
    16'h03e0: rd_data <= 32'h2703cb89;
    16'h03e1: rd_data <= 32'h2783fc04;
    16'h03e2: rd_data <= 32'h8f1dfcc4;
    16'h03e3: rd_data <= 32'heb842783;
    16'h03e4: rd_data <= 32'h2703c398;
    16'h03e5: rd_data <= 32'h2783fc44;
    16'h03e6: rd_data <= 32'h07b3fd04;
    16'h03e7: rd_data <= 32'h853e40f7;
    16'h03e8: rd_data <= 32'h14c12083;
    16'h03e9: rd_data <= 32'h14812403;
    16'h03ea: rd_data <= 32'h80826171;
    16'h03eb: rd_data <= 32'hd6067179;
    16'h03ec: rd_data <= 32'h1800d422;
    16'h03ed: rd_data <= 32'hfc042a23;
    16'h03ee: rd_data <= 32'h851367c5;
    16'h03ef: rd_data <= 32'hf0ef6d87;
    16'h03f0: rd_data <= 32'h07b7ce0f;
    16'h03f1: rd_data <= 32'h43940200;
    16'h03f2: rd_data <= 32'h020007b7;
    16'h03f3: rd_data <= 32'hff900737;
    16'h03f4: rd_data <= 32'h8f75177d;
    16'h03f5: rd_data <= 32'h67c5c398;
    16'h03f6: rd_data <= 32'h6e878513;
    16'h03f7: rd_data <= 32'hcc2ff0ef;
    16'h03f8: rd_data <= 32'hfd440793;
    16'h03f9: rd_data <= 32'h450185be;
    16'h03fa: rd_data <= 32'h87aa33c5;
    16'h03fb: rd_data <= 32'h853e45a1;
    16'h03fc: rd_data <= 32'hce4ff0ef;
    16'h03fd: rd_data <= 32'hf0ef4529;
    16'h03fe: rd_data <= 32'h47a1c76f;
    16'h03ff: rd_data <= 32'hfef42623;
    16'h0400: rd_data <= 32'h67c5a8a5;
    16'h0401: rd_data <= 32'h6ec78513;
    16'h0402: rd_data <= 32'hc96ff0ef;
    16'h0403: rd_data <= 32'hfec42783;
    16'h0404: rd_data <= 32'hf0ef853e;
    16'h0405: rd_data <= 32'h67c5d44f;
    16'h0406: rd_data <= 32'h6f478513;
    16'h0407: rd_data <= 32'hc82ff0ef;
    16'h0408: rd_data <= 32'hfec42783;
    16'h0409: rd_data <= 32'h0ff7f793;
    16'h040a: rd_data <= 32'hf0ef853e;
    16'h040b: rd_data <= 32'h07b7b0ef;
    16'h040c: rd_data <= 32'h43980200;
    16'h040d: rd_data <= 32'hff9007b7;
    16'h040e: rd_data <= 32'h76b317fd;
    16'h040f: rd_data <= 32'h07b700f7;
    16'h0410: rd_data <= 32'h07370200;
    16'h0411: rd_data <= 32'h8f550040;
    16'h0412: rd_data <= 32'h67c5c398;
    16'h0413: rd_data <= 32'h6e878513;
    16'h0414: rd_data <= 32'hc4eff0ef;
    16'h0415: rd_data <= 32'hfd440793;
    16'h0416: rd_data <= 32'h450185be;
    16'h0417: rd_data <= 32'h87aa33b5;
    16'h0418: rd_data <= 32'h853e45a1;
    16'h0419: rd_data <= 32'hc70ff0ef;
    16'h041a: rd_data <= 32'hf0ef4529;
    16'h041b: rd_data <= 32'h2783c02f;
    16'h041c: rd_data <= 32'h17fdfec4;
    16'h041d: rd_data <= 32'hfef42623;
    16'h041e: rd_data <= 32'hfec42783;
    16'h041f: rd_data <= 32'hf8f043e3;
    16'h0420: rd_data <= 32'h242347a1;
    16'h0421: rd_data <= 32'ha8a5fef4;
    16'h0422: rd_data <= 32'h851367c5;
    16'h0423: rd_data <= 32'hf0ef7007;
    16'h0424: rd_data <= 32'h2783c10f;
    16'h0425: rd_data <= 32'h853efe84;
    16'h0426: rd_data <= 32'hcbeff0ef;
    16'h0427: rd_data <= 32'h851367c5;
    16'h0428: rd_data <= 32'hf0ef70c7;
    16'h0429: rd_data <= 32'h2783bfcf;
    16'h042a: rd_data <= 32'hf793fe84;
    16'h042b: rd_data <= 32'h853e0ff7;
    16'h042c: rd_data <= 32'ha88ff0ef;
    16'h042d: rd_data <= 32'h020007b7;
    16'h042e: rd_data <= 32'h07b74398;
    16'h042f: rd_data <= 32'h17fdff90;
    16'h0430: rd_data <= 32'h00f776b3;
    16'h0431: rd_data <= 32'h020007b7;
    16'h0432: rd_data <= 32'h00500737;
    16'h0433: rd_data <= 32'hc3988f55;
    16'h0434: rd_data <= 32'h851367c5;
    16'h0435: rd_data <= 32'hf0ef6e87;
    16'h0436: rd_data <= 32'h0793bc8f;
    16'h0437: rd_data <= 32'h85befd44;
    16'h0438: rd_data <= 32'h31dd4501;
    16'h0439: rd_data <= 32'h45a187aa;
    16'h043a: rd_data <= 32'hf0ef853e;
    16'h043b: rd_data <= 32'h4529beaf;
    16'h043c: rd_data <= 32'hb7cff0ef;
    16'h043d: rd_data <= 32'hfe842783;
    16'h043e: rd_data <= 32'h242317fd;
    16'h043f: rd_data <= 32'h2783fef4;
    16'h0440: rd_data <= 32'h43e3fe84;
    16'h0441: rd_data <= 32'h47a1f8f0;
    16'h0442: rd_data <= 32'hfef42223;
    16'h0443: rd_data <= 32'h67c5a8a5;
    16'h0444: rd_data <= 32'h71478513;
    16'h0445: rd_data <= 32'hb8aff0ef;
    16'h0446: rd_data <= 32'hfe442783;
    16'h0447: rd_data <= 32'hf0ef853e;
    16'h0448: rd_data <= 32'h67c5c38f;
    16'h0449: rd_data <= 32'h6f478513;
    16'h044a: rd_data <= 32'hb76ff0ef;
    16'h044b: rd_data <= 32'hfe442783;
    16'h044c: rd_data <= 32'h0ff7f793;
    16'h044d: rd_data <= 32'hf0ef853e;
    16'h044e: rd_data <= 32'h07b7a02f;
    16'h044f: rd_data <= 32'h43980200;
    16'h0450: rd_data <= 32'hff9007b7;
    16'h0451: rd_data <= 32'h76b317fd;
    16'h0452: rd_data <= 32'h07b700f7;
    16'h0453: rd_data <= 32'h07370200;
    16'h0454: rd_data <= 32'h8f550020;
    16'h0455: rd_data <= 32'h67c5c398;
    16'h0456: rd_data <= 32'h6e878513;
    16'h0457: rd_data <= 32'hb42ff0ef;
    16'h0458: rd_data <= 32'hfd440793;
    16'h0459: rd_data <= 32'h450185be;
    16'h045a: rd_data <= 32'h87aa3185;
    16'h045b: rd_data <= 32'h853e45a1;
    16'h045c: rd_data <= 32'hb64ff0ef;
    16'h045d: rd_data <= 32'hf0ef4529;
    16'h045e: rd_data <= 32'h2783af6f;
    16'h045f: rd_data <= 32'h17fdfe44;
    16'h0460: rd_data <= 32'hfef42223;
    16'h0461: rd_data <= 32'hfe442783;
    16'h0462: rd_data <= 32'hf8f043e3;
    16'h0463: rd_data <= 32'h202347a1;
    16'h0464: rd_data <= 32'ha8a5fef4;
    16'h0465: rd_data <= 32'h851367c5;
    16'h0466: rd_data <= 32'hf0ef71c7;
    16'h0467: rd_data <= 32'h2783b04f;
    16'h0468: rd_data <= 32'h853efe04;
    16'h0469: rd_data <= 32'hbb2ff0ef;
    16'h046a: rd_data <= 32'h851367c5;
    16'h046b: rd_data <= 32'hf0ef70c7;
    16'h046c: rd_data <= 32'h2783af0f;
    16'h046d: rd_data <= 32'hf793fe04;
    16'h046e: rd_data <= 32'h853e0ff7;
    16'h046f: rd_data <= 32'h97cff0ef;
    16'h0470: rd_data <= 32'h020007b7;
    16'h0471: rd_data <= 32'h07b74398;
    16'h0472: rd_data <= 32'h17fdff90;
    16'h0473: rd_data <= 32'h00f776b3;
    16'h0474: rd_data <= 32'h020007b7;
    16'h0475: rd_data <= 32'h00300737;
    16'h0476: rd_data <= 32'hc3988f55;
    16'h0477: rd_data <= 32'h851367c5;
    16'h0478: rd_data <= 32'hf0ef6e87;
    16'h0479: rd_data <= 32'h0793abcf;
    16'h047a: rd_data <= 32'h85befd44;
    16'h047b: rd_data <= 32'h3ee94501;
    16'h047c: rd_data <= 32'h45a187aa;
    16'h047d: rd_data <= 32'hf0ef853e;
    16'h047e: rd_data <= 32'h4529adef;
    16'h047f: rd_data <= 32'ha70ff0ef;
    16'h0480: rd_data <= 32'hfe042783;
    16'h0481: rd_data <= 32'h202317fd;
    16'h0482: rd_data <= 32'h2783fef4;
    16'h0483: rd_data <= 32'h43e3fe04;
    16'h0484: rd_data <= 32'h47a1f8f0;
    16'h0485: rd_data <= 32'hfcf42e23;
    16'h0486: rd_data <= 32'h67c5a8a5;
    16'h0487: rd_data <= 32'h72878513;
    16'h0488: rd_data <= 32'ha7eff0ef;
    16'h0489: rd_data <= 32'hfdc42783;
    16'h048a: rd_data <= 32'hf0ef853e;
    16'h048b: rd_data <= 32'h67c5b2cf;
    16'h048c: rd_data <= 32'h70c78513;
    16'h048d: rd_data <= 32'ha6aff0ef;
    16'h048e: rd_data <= 32'hfdc42783;
    16'h048f: rd_data <= 32'h0ff7f793;
    16'h0490: rd_data <= 32'hf0ef853e;
    16'h0491: rd_data <= 32'h07b78f6f;
    16'h0492: rd_data <= 32'h43980200;
    16'h0493: rd_data <= 32'hff9007b7;
    16'h0494: rd_data <= 32'h76b317fd;
    16'h0495: rd_data <= 32'h07b700f7;
    16'h0496: rd_data <= 32'h07370200;
    16'h0497: rd_data <= 32'h8f550060;
    16'h0498: rd_data <= 32'h67c5c398;
    16'h0499: rd_data <= 32'h6e878513;
    16'h049a: rd_data <= 32'ha36ff0ef;
    16'h049b: rd_data <= 32'hfd440793;
    16'h049c: rd_data <= 32'h450185be;
    16'h049d: rd_data <= 32'h87aa3e91;
    16'h049e: rd_data <= 32'h853e45a1;
    16'h049f: rd_data <= 32'ha58ff0ef;
    16'h04a0: rd_data <= 32'hf0ef4529;
    16'h04a1: rd_data <= 32'h27839eaf;
    16'h04a2: rd_data <= 32'h17fdfdc4;
    16'h04a3: rd_data <= 32'hfcf42e23;
    16'h04a4: rd_data <= 32'hfdc42783;
    16'h04a5: rd_data <= 32'hf8f043e3;
    16'h04a6: rd_data <= 32'h2c2347a1;
    16'h04a7: rd_data <= 32'ha0bdfcf4;
    16'h04a8: rd_data <= 32'h851367c5;
    16'h04a9: rd_data <= 32'hf0ef7347;
    16'h04aa: rd_data <= 32'h27839f8f;
    16'h04ab: rd_data <= 32'h853efd84;
    16'h04ac: rd_data <= 32'haa6ff0ef;
    16'h04ad: rd_data <= 32'h851367c5;
    16'h04ae: rd_data <= 32'hf0ef67c7;
    16'h04af: rd_data <= 32'h27839e4f;
    16'h04b0: rd_data <= 32'hf793fd84;
    16'h04b1: rd_data <= 32'h853e0ff7;
    16'h04b2: rd_data <= 32'h870ff0ef;
    16'h04b3: rd_data <= 32'h020007b7;
    16'h04b4: rd_data <= 32'h07b74394;
    16'h04b5: rd_data <= 32'h07370200;
    16'h04b6: rd_data <= 32'h8f550070;
    16'h04b7: rd_data <= 32'h67c5c398;
    16'h04b8: rd_data <= 32'h6e878513;
    16'h04b9: rd_data <= 32'h9baff0ef;
    16'h04ba: rd_data <= 32'hfd440793;
    16'h04bb: rd_data <= 32'h450185be;
    16'h04bc: rd_data <= 32'h87aa3ce1;
    16'h04bd: rd_data <= 32'h853e45a1;
    16'h04be: rd_data <= 32'h9dcff0ef;
    16'h04bf: rd_data <= 32'hf0ef4529;
    16'h04c0: rd_data <= 32'h278396ef;
    16'h04c1: rd_data <= 32'h17fdfd84;
    16'h04c2: rd_data <= 32'hfcf42c23;
    16'h04c3: rd_data <= 32'hfd842783;
    16'h04c4: rd_data <= 32'hf8f048e3;
    16'h04c5: rd_data <= 32'h851367c5;
    16'h04c6: rd_data <= 32'hf0ef7447;
    16'h04c7: rd_data <= 32'h2783984f;
    16'h04c8: rd_data <= 32'h45a1fd44;
    16'h04c9: rd_data <= 32'hf0ef853e;
    16'h04ca: rd_data <= 32'h45299aef;
    16'h04cb: rd_data <= 32'h940ff0ef;
    16'h04cc: rd_data <= 32'h50b20001;
    16'h04cd: rd_data <= 32'h61455422;
    16'h04ce: rd_data <= 32'h11018082;
    16'h04cf: rd_data <= 32'hcc22ce06;
    16'h04d0: rd_data <= 32'h67c51000;
    16'h04d1: rd_data <= 32'h75878513;
    16'h04d2: rd_data <= 32'h956ff0ef;
    16'h04d3: rd_data <= 32'h4783a031;
    16'h04d4: rd_data <= 32'h853efef4;
    16'h04d5: rd_data <= 32'h918ff0ef;
    16'h04d6: rd_data <= 32'he02ff0ef;
    16'h04d7: rd_data <= 32'h07a387aa;
    16'h04d8: rd_data <= 32'h4703fef4;
    16'h04d9: rd_data <= 32'h0793fef4;
    16'h04da: rd_data <= 32'h12e30210;
    16'h04db: rd_data <= 32'h0001fef7;
    16'h04dc: rd_data <= 32'h446240f2;
    16'h04dd: rd_data <= 32'h80826105;
    16'h04de: rd_data <= 32'hce061101;
    16'h04df: rd_data <= 32'h1000cc22;
    16'h04e0: rd_data <= 32'h030007b7;
    16'h04e1: rd_data <= 32'hc398477d;
    16'h04e2: rd_data <= 32'h020007b7;
    16'h04e3: rd_data <= 32'h07130791;
    16'h04e4: rd_data <= 32'hc3980680;
    16'h04e5: rd_data <= 32'h851367c5;
    16'h04e6: rd_data <= 32'hf0ef7787;
    16'h04e7: rd_data <= 32'h07b7904f;
    16'h04e8: rd_data <= 32'h07130300;
    16'h04e9: rd_data <= 32'hc39803f0;
    16'h04ea: rd_data <= 32'heddfe0ef;
    16'h04eb: rd_data <= 32'h030007b7;
    16'h04ec: rd_data <= 32'h07f00713;
    16'h04ed: rd_data <= 32'h0001c398;
    16'h04ee: rd_data <= 32'h851367c5;
    16'h04ef: rd_data <= 32'hf0ef7847;
    16'h04f0: rd_data <= 32'h87aacf0f;
    16'h04f1: rd_data <= 32'h47b5873e;
    16'h04f2: rd_data <= 32'hfef718e3;
    16'h04f3: rd_data <= 32'h851367c5;
    16'h04f4: rd_data <= 32'hf0ef5fc7;
    16'h04f5: rd_data <= 32'h67c58ccf;
    16'h04f6: rd_data <= 32'h7a078513;
    16'h04f7: rd_data <= 32'h8c2ff0ef;
    16'h04f8: rd_data <= 32'h851367c5;
    16'h04f9: rd_data <= 32'hf0ef7c87;
    16'h04fa: rd_data <= 32'h67c58b8f;
    16'h04fb: rd_data <= 32'h7f078513;
    16'h04fc: rd_data <= 32'h8aeff0ef;
    16'h04fd: rd_data <= 32'h851367c9;
    16'h04fe: rd_data <= 32'hf0ef8147;
    16'h04ff: rd_data <= 32'h67c98a4f;
    16'h0500: rd_data <= 32'h83c78513;
    16'h0501: rd_data <= 32'h89aff0ef;
    16'h0502: rd_data <= 32'h851367c5;
    16'h0503: rd_data <= 32'hf0ef5fc7;
    16'h0504: rd_data <= 32'h67c9890f;
    16'h0505: rd_data <= 32'h86478513;
    16'h0506: rd_data <= 32'h886ff0ef;
    16'h0507: rd_data <= 32'h08000513;
    16'h0508: rd_data <= 32'h936ff0ef;
    16'h0509: rd_data <= 32'h851367c9;
    16'h050a: rd_data <= 32'hf0ef8747;
    16'h050b: rd_data <= 32'h67c5874f;
    16'h050c: rd_data <= 32'h5fc78513;
    16'h050d: rd_data <= 32'h86aff0ef;
    16'h050e: rd_data <= 32'he44ff0ef;
    16'h050f: rd_data <= 32'h851367c5;
    16'h0510: rd_data <= 32'hf0ef5fc7;
    16'h0511: rd_data <= 32'hf0ef85cf;
    16'h0512: rd_data <= 32'h67c5d2cf;
    16'h0513: rd_data <= 32'h5fc78513;
    16'h0514: rd_data <= 32'h84eff0ef;
    16'h0515: rd_data <= 32'h851367c5;
    16'h0516: rd_data <= 32'hf0ef5fc7;
    16'h0517: rd_data <= 32'h67c9844f;
    16'h0518: rd_data <= 32'h87c78513;
    16'h0519: rd_data <= 32'h83aff0ef;
    16'h051a: rd_data <= 32'h851367c5;
    16'h051b: rd_data <= 32'hf0ef5fc7;
    16'h051c: rd_data <= 32'h67c9830f;
    16'h051d: rd_data <= 32'h89078513;
    16'h051e: rd_data <= 32'h826ff0ef;
    16'h051f: rd_data <= 32'h851367c9;
    16'h0520: rd_data <= 32'hf0ef8ac7;
    16'h0521: rd_data <= 32'h67c981cf;
    16'h0522: rd_data <= 32'h8cc78513;
    16'h0523: rd_data <= 32'h812ff0ef;
    16'h0524: rd_data <= 32'h851367c9;
    16'h0525: rd_data <= 32'hf0ef8ec7;
    16'h0526: rd_data <= 32'h67c9808f;
    16'h0527: rd_data <= 32'h90c78513;
    16'h0528: rd_data <= 32'hffffe0ef;
    16'h0529: rd_data <= 32'h851367c9;
    16'h052a: rd_data <= 32'he0ef92c7;
    16'h052b: rd_data <= 32'h67c9ff5f;
    16'h052c: rd_data <= 32'h94c78513;
    16'h052d: rd_data <= 32'hfebfe0ef;
    16'h052e: rd_data <= 32'h851367c9;
    16'h052f: rd_data <= 32'he0ef9707;
    16'h0530: rd_data <= 32'h67c9fe1f;
    16'h0531: rd_data <= 32'h99478513;
    16'h0532: rd_data <= 32'hfd7fe0ef;
    16'h0533: rd_data <= 32'h851367c9;
    16'h0534: rd_data <= 32'he0ef9b47;
    16'h0535: rd_data <= 32'h67c9fcdf;
    16'h0536: rd_data <= 32'h9c878513;
    16'h0537: rd_data <= 32'hfc3fe0ef;
    16'h0538: rd_data <= 32'h851367c9;
    16'h0539: rd_data <= 32'he0ef9e07;
    16'h053a: rd_data <= 32'h67c5fb9f;
    16'h053b: rd_data <= 32'h5fc78513;
    16'h053c: rd_data <= 32'hfaffe0ef;
    16'h053d: rd_data <= 32'h262347a9;
    16'h053e: rd_data <= 32'ha0d1fef4;
    16'h053f: rd_data <= 32'h851367c9;
    16'h0540: rd_data <= 32'he0ef9f47;
    16'h0541: rd_data <= 32'hf0eff9df;
    16'h0542: rd_data <= 32'h87aac54f;
    16'h0543: rd_data <= 32'hfef405a3;
    16'h0544: rd_data <= 32'hfeb44703;
    16'h0545: rd_data <= 32'h02000793;
    16'h0546: rd_data <= 32'h00e7fd63;
    16'h0547: rd_data <= 32'hfeb44703;
    16'h0548: rd_data <= 32'h07e00793;
    16'h0549: rd_data <= 32'h00e7e763;
    16'h054a: rd_data <= 32'hfeb44783;
    16'h054b: rd_data <= 32'he0ef853e;
    16'h054c: rd_data <= 32'h67c5f3ff;
    16'h054d: rd_data <= 32'h5fc78513;
    16'h054e: rd_data <= 32'hf67fe0ef;
    16'h054f: rd_data <= 32'hfeb44783;
    16'h0550: rd_data <= 32'hfd078793;
    16'h0551: rd_data <= 32'h03500713;
    16'h0552: rd_data <= 32'h06f76463;
    16'h0553: rd_data <= 32'h00279713;
    16'h0554: rd_data <= 32'h879367c9;
    16'h0555: rd_data <= 32'h97baa007;
    16'h0556: rd_data <= 32'h8782439c;
    16'h0557: rd_data <= 32'hea8ff0ef;
    16'h0558: rd_data <= 32'hf0efa8b1;
    16'h0559: rd_data <= 32'ha899fcaf;
    16'h055a: rd_data <= 32'he65fe0ef;
    16'h055b: rd_data <= 32'he0efa881;
    16'h055c: rd_data <= 32'ha0a9e81f;
    16'h055d: rd_data <= 32'hea5fe0ef;
    16'h055e: rd_data <= 32'he0efa091;
    16'h055f: rd_data <= 32'ha83dec9f;
    16'h0560: rd_data <= 32'h020007b7;
    16'h0561: rd_data <= 32'h07b74394;
    16'h0562: rd_data <= 32'h07370200;
    16'h0563: rd_data <= 32'h8f350010;
    16'h0564: rd_data <= 32'ha02dc398;
    16'h0565: rd_data <= 32'h45054581;
    16'h0566: rd_data <= 32'ha00d3805;
    16'h0567: rd_data <= 32'ha8393c01;
    16'h0568: rd_data <= 32'hcdcff0ef;
    16'h0569: rd_data <= 32'hf0efa821;
    16'h056a: rd_data <= 32'ha809bccf;
    16'h056b: rd_data <= 32'ha0393379;
    16'h056c: rd_data <= 32'hfec42783;
    16'h056d: rd_data <= 32'h262317fd;
    16'h056e: rd_data <= 32'ha011fef4;
    16'h056f: rd_data <= 32'h2783a029;
    16'h0570: rd_data <= 32'h4de3fec4;
    16'h0571: rd_data <= 32'hb579f2f0;
    16'h0572: rd_data <= 32'h33323130;
    16'h0573: rd_data <= 32'h37363534;
    16'h0574: rd_data <= 32'h62613938;
    16'h0575: rd_data <= 32'h66656463;
    16'h0576: rd_data <= 32'h00000000;
    16'h0577: rd_data <= 32'h30313d3e;
    16'h0578: rd_data <= 32'h00003030;
    16'h0579: rd_data <= 32'h20495053;
    16'h057a: rd_data <= 32'h74617453;
    16'h057b: rd_data <= 32'h000a3a65;
    16'h057c: rd_data <= 32'h414c2020;
    16'h057d: rd_data <= 32'h434e4554;
    16'h057e: rd_data <= 32'h00002059;
    16'h057f: rd_data <= 32'h0000000a;
    16'h0580: rd_data <= 32'h44442020;
    16'h0581: rd_data <= 32'h00002052;
    16'h0582: rd_data <= 32'h000a4e4f;
    16'h0583: rd_data <= 32'h0a46464f;
    16'h0584: rd_data <= 32'h00000000;
    16'h0585: rd_data <= 32'h53512020;
    16'h0586: rd_data <= 32'h00204950;
    16'h0587: rd_data <= 32'h52432020;
    16'h0588: rd_data <= 32'h0000204d;
    16'h0589: rd_data <= 32'h6e6e7552;
    16'h058a: rd_data <= 32'h20676e69;
    16'h058b: rd_data <= 32'h746d656d;
    16'h058c: rd_data <= 32'h20747365;
    16'h058d: rd_data <= 32'h00000000;
    16'h058e: rd_data <= 32'h2a2a2a20;
    16'h058f: rd_data <= 32'h4c494146;
    16'h0590: rd_data <= 32'h57204445;
    16'h0591: rd_data <= 32'h2a44524f;
    16'h0592: rd_data <= 32'h61202a2a;
    16'h0593: rd_data <= 32'h00002074;
    16'h0594: rd_data <= 32'h0000002e;
    16'h0595: rd_data <= 32'h2a2a2a20;
    16'h0596: rd_data <= 32'h4c494146;
    16'h0597: rd_data <= 32'h42204445;
    16'h0598: rd_data <= 32'h2a455459;
    16'h0599: rd_data <= 32'h61202a2a;
    16'h059a: rd_data <= 32'h00002074;
    16'h059b: rd_data <= 32'h73617020;
    16'h059c: rd_data <= 32'h0a646573;
    16'h059d: rd_data <= 32'h00000000;
    16'h059e: rd_data <= 32'h00007830;
    16'h059f: rd_data <= 32'h00000020;
    16'h05a0: rd_data <= 32'h00783020;
    16'h05a1: rd_data <= 32'h56315253;
    16'h05a2: rd_data <= 32'h00000000;
    16'h05a3: rd_data <= 32'h56325253;
    16'h05a4: rd_data <= 32'h00000000;
    16'h05a5: rd_data <= 32'h56315243;
    16'h05a6: rd_data <= 32'h00000000;
    16'h05a7: rd_data <= 32'h56325243;
    16'h05a8: rd_data <= 32'h00000000;
    16'h05a9: rd_data <= 32'h56335243;
    16'h05aa: rd_data <= 32'h00000000;
    16'h05ab: rd_data <= 32'h504c4456;
    16'h05ac: rd_data <= 32'h00000000;
    16'h05ad: rd_data <= 32'h6c637943;
    16'h05ae: rd_data <= 32'h203a7365;
    16'h05af: rd_data <= 32'h00007830;
    16'h05b0: rd_data <= 32'h74736e49;
    16'h05b1: rd_data <= 32'h203a736e;
    16'h05b2: rd_data <= 32'h00007830;
    16'h05b3: rd_data <= 32'h736b6843;
    16'h05b4: rd_data <= 32'h203a6d75;
    16'h05b5: rd_data <= 32'h00007830;
    16'h05b6: rd_data <= 32'h61666564;
    16'h05b7: rd_data <= 32'h20746c75;
    16'h05b8: rd_data <= 32'h20202020;
    16'h05b9: rd_data <= 32'h00202020;
    16'h05ba: rd_data <= 32'h0000203a;
    16'h05bb: rd_data <= 32'h69707364;
    16'h05bc: rd_data <= 32'h0000002d;
    16'h05bd: rd_data <= 32'h20202020;
    16'h05be: rd_data <= 32'h20202020;
    16'h05bf: rd_data <= 32'h00000020;
    16'h05c0: rd_data <= 32'h69707364;
    16'h05c1: rd_data <= 32'h6d72632d;
    16'h05c2: rd_data <= 32'h0000002d;
    16'h05c3: rd_data <= 32'h20202020;
    16'h05c4: rd_data <= 32'h00000020;
    16'h05c5: rd_data <= 32'h69707371;
    16'h05c6: rd_data <= 32'h0000002d;
    16'h05c7: rd_data <= 32'h69707371;
    16'h05c8: rd_data <= 32'h6d72632d;
    16'h05c9: rd_data <= 32'h0000002d;
    16'h05ca: rd_data <= 32'h69707371;
    16'h05cb: rd_data <= 32'h7264642d;
    16'h05cc: rd_data <= 32'h0000002d;
    16'h05cd: rd_data <= 32'h69707371;
    16'h05ce: rd_data <= 32'h7264642d;
    16'h05cf: rd_data <= 32'h6d72632d;
    16'h05d0: rd_data <= 32'h0000002d;
    16'h05d1: rd_data <= 32'h74736e69;
    16'h05d2: rd_data <= 32'h2020736e;
    16'h05d3: rd_data <= 32'h20202020;
    16'h05d4: rd_data <= 32'h3a202020;
    16'h05d5: rd_data <= 32'h00000020;
    16'h05d6: rd_data <= 32'h75746552;
    16'h05d7: rd_data <= 32'h74206e72;
    16'h05d8: rd_data <= 32'h656d206f;
    16'h05d9: rd_data <= 32'h6220756e;
    16'h05da: rd_data <= 32'h65732079;
    16'h05db: rd_data <= 32'h6e69646e;
    16'h05dc: rd_data <= 32'h21272067;
    16'h05dd: rd_data <= 32'h000a0a27;
    16'h05de: rd_data <= 32'h746f6f42;
    16'h05df: rd_data <= 32'h2e676e69;
    16'h05e0: rd_data <= 32'h00000a2e;
    16'h05e1: rd_data <= 32'h73657250;
    16'h05e2: rd_data <= 32'h4e452073;
    16'h05e3: rd_data <= 32'h20524554;
    16'h05e4: rd_data <= 32'h63206f74;
    16'h05e5: rd_data <= 32'h69746e6f;
    16'h05e6: rd_data <= 32'h2e65756e;
    16'h05e7: rd_data <= 32'h00000a2e;
    16'h05e8: rd_data <= 32'h5f5f2020;
    16'h05e9: rd_data <= 32'h20205f5f;
    16'h05ea: rd_data <= 32'h2020205f;
    16'h05eb: rd_data <= 32'h20202020;
    16'h05ec: rd_data <= 32'h5f202020;
    16'h05ed: rd_data <= 32'h205f5f5f;
    16'h05ee: rd_data <= 32'h20202020;
    16'h05ef: rd_data <= 32'h20202020;
    16'h05f0: rd_data <= 32'h5f5f5f5f;
    16'h05f1: rd_data <= 32'h0000000a;
    16'h05f2: rd_data <= 32'h20207c20;
    16'h05f3: rd_data <= 32'h285c205f;
    16'h05f4: rd_data <= 32'h5f20295f;
    16'h05f5: rd_data <= 32'h5f205f5f;
    16'h05f6: rd_data <= 32'h202f5f5f;
    16'h05f7: rd_data <= 32'h7c5f5f5f;
    16'h05f8: rd_data <= 32'h5f5f2020;
    16'h05f9: rd_data <= 32'h2f20205f;
    16'h05fa: rd_data <= 32'h5f5f5f20;
    16'h05fb: rd_data <= 32'h00000a7c;
    16'h05fc: rd_data <= 32'h7c207c20;
    16'h05fd: rd_data <= 32'h7c20295f;
    16'h05fe: rd_data <= 32'h202f7c20;
    16'h05ff: rd_data <= 32'h202f5f5f;
    16'h0600: rd_data <= 32'h5f5c205f;
    16'h0601: rd_data <= 32'h5c205f5f;
    16'h0602: rd_data <= 32'h5f202f20;
    16'h0603: rd_data <= 32'h207c5c20;
    16'h0604: rd_data <= 32'h00000a7c;
    16'h0605: rd_data <= 32'h20207c20;
    16'h0606: rd_data <= 32'h7c2f5f5f;
    16'h0607: rd_data <= 32'h28207c20;
    16'h0608: rd_data <= 32'h28207c5f;
    16'h0609: rd_data <= 32'h7c20295f;
    16'h060a: rd_data <= 32'h20295f5f;
    16'h060b: rd_data <= 32'h5f28207c;
    16'h060c: rd_data <= 32'h207c2029;
    16'h060d: rd_data <= 32'h5f5f5f7c;
    16'h060e: rd_data <= 32'h0000000a;
    16'h060f: rd_data <= 32'h7c5f7c20;
    16'h0610: rd_data <= 32'h7c202020;
    16'h0611: rd_data <= 32'h5f5c7c5f;
    16'h0612: rd_data <= 32'h5f5c5f5f;
    16'h0613: rd_data <= 32'h5f2f5f5f;
    16'h0614: rd_data <= 32'h2f5f5f5f;
    16'h0615: rd_data <= 32'h5f5f5c20;
    16'h0616: rd_data <= 32'h5c202f5f;
    16'h0617: rd_data <= 32'h5f5f5f5f;
    16'h0618: rd_data <= 32'h00000a7c;
    16'h0619: rd_data <= 32'h61746f54;
    16'h061a: rd_data <= 32'h656d206c;
    16'h061b: rd_data <= 32'h79726f6d;
    16'h061c: rd_data <= 32'h0000203a;
    16'h061d: rd_data <= 32'h42694b20;
    16'h061e: rd_data <= 32'h0000000a;
    16'h061f: rd_data <= 32'h656c6553;
    16'h0620: rd_data <= 32'h61207463;
    16'h0621: rd_data <= 32'h6361206e;
    16'h0622: rd_data <= 32'h6e6f6974;
    16'h0623: rd_data <= 32'h00000a3a;
    16'h0624: rd_data <= 32'h5b202020;
    16'h0625: rd_data <= 32'h52205d31;
    16'h0626: rd_data <= 32'h20646165;
    16'h0627: rd_data <= 32'h20495053;
    16'h0628: rd_data <= 32'h73616c46;
    16'h0629: rd_data <= 32'h44492068;
    16'h062a: rd_data <= 32'h0000000a;
    16'h062b: rd_data <= 32'h5b202020;
    16'h062c: rd_data <= 32'h52205d32;
    16'h062d: rd_data <= 32'h20646165;
    16'h062e: rd_data <= 32'h20495053;
    16'h062f: rd_data <= 32'h666e6f43;
    16'h0630: rd_data <= 32'h52206769;
    16'h0631: rd_data <= 32'h0a736765;
    16'h0632: rd_data <= 32'h00000000;
    16'h0633: rd_data <= 32'h5b202020;
    16'h0634: rd_data <= 32'h53205d33;
    16'h0635: rd_data <= 32'h63746977;
    16'h0636: rd_data <= 32'h6f742068;
    16'h0637: rd_data <= 32'h66656420;
    16'h0638: rd_data <= 32'h746c7561;
    16'h0639: rd_data <= 32'h646f6d20;
    16'h063a: rd_data <= 32'h00000a65;
    16'h063b: rd_data <= 32'h5b202020;
    16'h063c: rd_data <= 32'h53205d34;
    16'h063d: rd_data <= 32'h63746977;
    16'h063e: rd_data <= 32'h6f742068;
    16'h063f: rd_data <= 32'h61754420;
    16'h0640: rd_data <= 32'h2f49206c;
    16'h0641: rd_data <= 32'h6f6d204f;
    16'h0642: rd_data <= 32'h000a6564;
    16'h0643: rd_data <= 32'h5b202020;
    16'h0644: rd_data <= 32'h53205d35;
    16'h0645: rd_data <= 32'h63746977;
    16'h0646: rd_data <= 32'h6f742068;
    16'h0647: rd_data <= 32'h61755120;
    16'h0648: rd_data <= 32'h2f492064;
    16'h0649: rd_data <= 32'h6f6d204f;
    16'h064a: rd_data <= 32'h000a6564;
    16'h064b: rd_data <= 32'h5b202020;
    16'h064c: rd_data <= 32'h53205d36;
    16'h064d: rd_data <= 32'h63746977;
    16'h064e: rd_data <= 32'h6f742068;
    16'h064f: rd_data <= 32'h61755120;
    16'h0650: rd_data <= 32'h44442064;
    16'h0651: rd_data <= 32'h6f6d2052;
    16'h0652: rd_data <= 32'h000a6564;
    16'h0653: rd_data <= 32'h5b202020;
    16'h0654: rd_data <= 32'h54205d37;
    16'h0655: rd_data <= 32'h6c67676f;
    16'h0656: rd_data <= 32'h6f632065;
    16'h0657: rd_data <= 32'h6e69746e;
    16'h0658: rd_data <= 32'h73756f75;
    16'h0659: rd_data <= 32'h61657220;
    16'h065a: rd_data <= 32'h6f6d2064;
    16'h065b: rd_data <= 32'h000a6564;
    16'h065c: rd_data <= 32'h5b202020;
    16'h065d: rd_data <= 32'h52205d39;
    16'h065e: rd_data <= 32'h73206e75;
    16'h065f: rd_data <= 32'h6c706d69;
    16'h0660: rd_data <= 32'h69747369;
    16'h0661: rd_data <= 32'h65622063;
    16'h0662: rd_data <= 32'h6d68636e;
    16'h0663: rd_data <= 32'h0a6b7261;
    16'h0664: rd_data <= 32'h00000000;
    16'h0665: rd_data <= 32'h5b202020;
    16'h0666: rd_data <= 32'h42205d30;
    16'h0667: rd_data <= 32'h68636e65;
    16'h0668: rd_data <= 32'h6b72616d;
    16'h0669: rd_data <= 32'h6c6c6120;
    16'h066a: rd_data <= 32'h6e6f6320;
    16'h066b: rd_data <= 32'h73676966;
    16'h066c: rd_data <= 32'h0000000a;
    16'h066d: rd_data <= 32'h5b202020;
    16'h066e: rd_data <= 32'h52205d4d;
    16'h066f: rd_data <= 32'h4d206e75;
    16'h0670: rd_data <= 32'h65746d65;
    16'h0671: rd_data <= 32'h000a7473;
    16'h0672: rd_data <= 32'h5b202020;
    16'h0673: rd_data <= 32'h50205d53;
    16'h0674: rd_data <= 32'h746e6972;
    16'h0675: rd_data <= 32'h49505320;
    16'h0676: rd_data <= 32'h61747320;
    16'h0677: rd_data <= 32'h000a6574;
    16'h0678: rd_data <= 32'h5b202020;
    16'h0679: rd_data <= 32'h45205d65;
    16'h067a: rd_data <= 32'h206f6863;
    16'h067b: rd_data <= 32'h54524155;
    16'h067c: rd_data <= 32'h0000000a;
    16'h067d: rd_data <= 32'h6d6d6f43;
    16'h067e: rd_data <= 32'h3e646e61;
    16'h067f: rd_data <= 32'h00000020;
    16'h0680: rd_data <= 32'h0001159c;
    16'h0681: rd_data <= 32'h0001155c;
    16'h0682: rd_data <= 32'h00011562;
    16'h0683: rd_data <= 32'h00011568;
    16'h0684: rd_data <= 32'h0001156e;
    16'h0685: rd_data <= 32'h00011574;
    16'h0686: rd_data <= 32'h0001157a;
    16'h0687: rd_data <= 32'h00011580;
    16'h0688: rd_data <= 32'h000115b0;
    16'h0689: rd_data <= 32'h00011594;
    16'h068a: rd_data <= 32'h000115b0;
    16'h068b: rd_data <= 32'h000115b0;
    16'h068c: rd_data <= 32'h000115b0;
    16'h068d: rd_data <= 32'h000115b0;
    16'h068e: rd_data <= 32'h000115b0;
    16'h068f: rd_data <= 32'h000115b0;
    16'h0690: rd_data <= 32'h000115b0;
    16'h0691: rd_data <= 32'h000115b0;
    16'h0692: rd_data <= 32'h000115b0;
    16'h0693: rd_data <= 32'h000115b0;
    16'h0694: rd_data <= 32'h000115b0;
    16'h0695: rd_data <= 32'h000115b0;
    16'h0696: rd_data <= 32'h000115b0;
    16'h0697: rd_data <= 32'h000115b0;
    16'h0698: rd_data <= 32'h000115b0;
    16'h0699: rd_data <= 32'h000115b0;
    16'h069a: rd_data <= 32'h000115b0;
    16'h069b: rd_data <= 32'h000115b0;
    16'h069c: rd_data <= 32'h000115b0;
    16'h069d: rd_data <= 32'h000115a0;
    16'h069e: rd_data <= 32'h000115b0;
    16'h069f: rd_data <= 32'h000115b0;
    16'h06a0: rd_data <= 32'h000115a6;
    16'h06a1: rd_data <= 32'h000115b0;
    16'h06a2: rd_data <= 32'h000115b0;
    16'h06a3: rd_data <= 32'h000115b0;
    16'h06a4: rd_data <= 32'h000115b0;
    16'h06a5: rd_data <= 32'h000115b0;
    16'h06a6: rd_data <= 32'h000115b0;
    16'h06a7: rd_data <= 32'h000115b0;
    16'h06a8: rd_data <= 32'h000115b0;
    16'h06a9: rd_data <= 32'h000115b0;
    16'h06aa: rd_data <= 32'h000115b0;
    16'h06ab: rd_data <= 32'h000115b0;
    16'h06ac: rd_data <= 32'h000115b0;
    16'h06ad: rd_data <= 32'h000115b0;
    16'h06ae: rd_data <= 32'h000115b0;
    16'h06af: rd_data <= 32'h000115b0;
    16'h06b0: rd_data <= 32'h000115b0;
    16'h06b1: rd_data <= 32'h000115b0;
    16'h06b2: rd_data <= 32'h000115b0;
    16'h06b3: rd_data <= 32'h000115b0;
    16'h06b4: rd_data <= 32'h000115b0;
    16'h06b5: rd_data <= 32'h000115ac;
    default: rd_data <= 32'h00000000;
  endcase

endmodule
